`define PI 3.14159265359
`define SCALE 1024

`define INT_RNS_DELTA_64 1968032985454108850
`define RNS_MIDDLE_POINT_64 8239355544127721383
`define MAX_NUM_64 16478711088255442766

`define A0 8239355544127721383
`define A1 2811533645389554216
`define A2 12636141686509778982
`define A3 3702265486788667758
`define A4 7483781454928236016
`define A5 636516737314587918
`define A6 6412218122208184842
`define A7 752140340127841786
`define A8 6762180247371755398

`define B0 2
`define B1 211
`define B2 223
`define B3 227
`define B4 229
`define B5 233
`define B6 239
`define B7 241
`define B8 251