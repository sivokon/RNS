`define INT_RNS_DELTA 926404979
`define RNS_MIDDLE_POINT 1684281159

`define B0 233
`define B1 239
`define B2 241
`define B3 251
