// this file is placeholder for common code
`define PI 3.14159265359
`define SCALE 1024
