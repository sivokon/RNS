// this file is placeholder for common code
`define PI 3.14159265359
`define SCALE 1024

`define INT_RNS_DELTA 926404979
`define RNS_MIDDLE_POINT 1684281159
